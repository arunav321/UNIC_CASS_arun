magic
tech sky130A
magscale 1 2
timestamp 1727354763
<< checkpaint >>
rect 1270 -3284 4212 94
<< error_s >>
rect 298 -865 333 -831
rect 299 -884 333 -865
rect 129 -933 187 -927
rect 129 -967 141 -933
rect 129 -973 187 -967
rect 101 -1001 200 -1000
rect 318 -1617 333 -884
rect 352 -918 387 -884
rect 667 -918 702 -884
rect 352 -1617 386 -918
rect 668 -937 702 -918
rect 498 -986 556 -980
rect 498 -1020 510 -986
rect 498 -1026 556 -1020
rect 498 -1534 556 -1528
rect 498 -1568 510 -1534
rect 498 -1574 556 -1568
rect 352 -1651 367 -1617
rect 687 -1670 702 -937
rect 721 -971 756 -937
rect 1036 -971 1071 -937
rect 721 -1670 755 -971
rect 1037 -990 1071 -971
rect 867 -1039 925 -1033
rect 867 -1073 879 -1039
rect 867 -1079 925 -1073
rect 867 -1587 925 -1581
rect 867 -1621 879 -1587
rect 867 -1627 925 -1621
rect 721 -1704 736 -1670
rect 1056 -1723 1071 -990
rect 1090 -1024 1125 -990
rect 1405 -1024 1440 -990
rect 1090 -1723 1124 -1024
rect 1406 -1043 1440 -1024
rect 1236 -1092 1294 -1086
rect 1236 -1126 1248 -1092
rect 1236 -1132 1294 -1126
rect 1236 -1640 1294 -1634
rect 1236 -1674 1248 -1640
rect 1236 -1680 1294 -1674
rect 1090 -1757 1105 -1723
rect 1425 -1776 1440 -1043
rect 1459 -1077 1494 -1043
rect 1774 -1077 1809 -1043
rect 1459 -1776 1493 -1077
rect 1775 -1096 1809 -1077
rect 1605 -1145 1663 -1139
rect 1605 -1179 1617 -1145
rect 1605 -1185 1663 -1179
rect 1605 -1693 1663 -1687
rect 1605 -1727 1617 -1693
rect 1605 -1733 1663 -1727
rect 1459 -1810 1474 -1776
rect 1794 -1829 1809 -1096
rect 1828 -1130 1863 -1096
rect 2143 -1130 2178 -1096
rect 1828 -1829 1862 -1130
rect 2144 -1149 2178 -1130
rect 1974 -1198 2032 -1192
rect 1974 -1232 1986 -1198
rect 1974 -1238 2032 -1232
rect 1974 -1746 2032 -1740
rect 1974 -1780 1986 -1746
rect 1974 -1786 2032 -1780
rect 1828 -1863 1843 -1829
rect 2163 -1882 2178 -1149
rect 2197 -1183 2232 -1149
rect 2512 -1183 2547 -1149
rect 2197 -1882 2231 -1183
rect 2513 -1202 2547 -1183
rect 2343 -1251 2401 -1245
rect 2343 -1285 2355 -1251
rect 2343 -1291 2401 -1285
rect 2343 -1799 2401 -1793
rect 2343 -1833 2355 -1799
rect 2343 -1839 2401 -1833
rect 2197 -1916 2212 -1882
rect 2532 -1935 2547 -1202
rect 2566 -1236 2601 -1202
rect 2881 -1236 2916 -1219
rect 2566 -1935 2600 -1236
rect 2882 -1237 2916 -1236
rect 2882 -1273 2952 -1237
rect 2712 -1304 2770 -1298
rect 2712 -1338 2724 -1304
rect 2899 -1307 2970 -1273
rect 3250 -1307 3285 -1273
rect 2712 -1344 2770 -1338
rect 2712 -1852 2770 -1846
rect 2712 -1886 2724 -1852
rect 2712 -1892 2770 -1886
rect 2566 -1969 2581 -1935
rect 2899 -1988 2969 -1307
rect 3251 -1326 3285 -1307
rect 3081 -1375 3139 -1369
rect 3081 -1409 3093 -1375
rect 3081 -1415 3139 -1409
rect 3081 -1905 3139 -1899
rect 3081 -1939 3093 -1905
rect 3081 -1945 3139 -1939
rect 2899 -2024 2952 -1988
rect 3270 -2041 3285 -1326
rect 3304 -1360 3339 -1326
rect 3619 -1360 3654 -1326
rect 3304 -2041 3338 -1360
rect 3620 -1379 3654 -1360
rect 3450 -1428 3508 -1422
rect 3450 -1462 3462 -1428
rect 3450 -1468 3508 -1462
rect 3450 -1958 3508 -1952
rect 3450 -1992 3462 -1958
rect 3450 -1998 3508 -1992
rect 3304 -2075 3319 -2041
rect 3639 -2094 3654 -1379
rect 3673 -1413 3708 -1379
rect 3988 -1413 4023 -1379
rect 3673 -2094 3707 -1413
rect 3989 -1432 4023 -1413
rect 3819 -1481 3877 -1475
rect 3819 -1515 3831 -1481
rect 3819 -1521 3877 -1515
rect 3819 -2011 3877 -2005
rect 3819 -2045 3831 -2011
rect 3819 -2051 3877 -2045
rect 3673 -2128 3688 -2094
rect 4008 -2147 4023 -1432
rect 4042 -1466 4077 -1432
rect 4357 -1466 4392 -1432
rect 4042 -2147 4076 -1466
rect 4358 -1485 4392 -1466
rect 4188 -1534 4246 -1528
rect 4188 -1568 4200 -1534
rect 4188 -1574 4246 -1568
rect 4188 -2064 4246 -2058
rect 4188 -2098 4200 -2064
rect 4188 -2104 4246 -2098
rect 4042 -2181 4057 -2147
rect 4377 -2200 4392 -1485
rect 4411 -1519 4446 -1485
rect 4726 -1519 4761 -1485
rect 4411 -2200 4445 -1519
rect 4727 -1538 4761 -1519
rect 4557 -1587 4615 -1581
rect 4557 -1621 4569 -1587
rect 4557 -1627 4615 -1621
rect 4557 -2117 4615 -2111
rect 4557 -2151 4569 -2117
rect 4557 -2157 4615 -2151
rect 4411 -2234 4426 -2200
rect 4746 -2253 4761 -1538
rect 4780 -1572 4815 -1538
rect 5095 -1572 5130 -1538
rect 4780 -2253 4814 -1572
rect 5096 -1591 5130 -1572
rect 4926 -1640 4984 -1634
rect 4926 -1674 4938 -1640
rect 4926 -1680 4984 -1674
rect 4926 -2170 4984 -2164
rect 4926 -2204 4938 -2170
rect 4926 -2210 4984 -2204
rect 4780 -2287 4795 -2253
rect 5115 -2306 5130 -1591
rect 5149 -1625 5184 -1591
rect 5464 -1625 5499 -1591
rect 5149 -2306 5183 -1625
rect 5465 -1644 5499 -1625
rect 5295 -1693 5353 -1687
rect 5295 -1727 5307 -1693
rect 5295 -1733 5353 -1727
rect 5295 -2223 5353 -2217
rect 5295 -2257 5307 -2223
rect 5295 -2263 5353 -2257
rect 5149 -2340 5164 -2306
rect 5484 -2359 5499 -1644
rect 5518 -1678 5553 -1644
rect 5833 -1678 5868 -1644
rect 5518 -2359 5552 -1678
rect 5834 -1697 5868 -1678
rect 5664 -1746 5722 -1740
rect 5664 -1780 5676 -1746
rect 5664 -1786 5722 -1780
rect 5664 -2276 5722 -2270
rect 5664 -2310 5676 -2276
rect 5664 -2316 5722 -2310
rect 5518 -2393 5533 -2359
rect 5853 -2412 5868 -1697
rect 5887 -1731 5922 -1697
rect 6202 -1731 6237 -1697
rect 5887 -2412 5921 -1731
rect 6203 -1750 6237 -1731
rect 6033 -1799 6091 -1793
rect 6033 -1833 6045 -1799
rect 6033 -1839 6091 -1833
rect 6033 -2329 6091 -2323
rect 6033 -2363 6045 -2329
rect 6033 -2369 6091 -2363
rect 5887 -2446 5902 -2412
rect 6222 -2465 6237 -1750
rect 6256 -1784 6291 -1750
rect 6256 -2465 6290 -1784
rect 6402 -1852 6460 -1846
rect 6402 -1886 6414 -1852
rect 6402 -1892 6460 -1886
rect 6402 -2382 6460 -2376
rect 6402 -2416 6414 -2382
rect 6402 -2422 6460 -2416
rect 6256 -2499 6271 -2465
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__pfet_01v8_WGVR8J  X0
timestamp 0
transform 1 0 2372 0 1 -1542
box -211 -429 211 429
use sky130_fd_pr__pfet_01v8_6FCS7L  X2
timestamp 0
transform 1 0 896 0 1 -1330
box -211 -429 211 429
use sky130_fd_pr__pfet_01v8_ETRZ5W  X3
timestamp 0
transform 1 0 1265 0 1 -1383
box -211 -429 211 429
use sky130_fd_pr__nfet_01v8_GBWJGK  X4
timestamp 0
transform 1 0 5324 0 1 -1975
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X5
timestamp 0
transform 1 0 5693 0 1 -2028
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_UJAU4L  X6
timestamp 0
transform 1 0 6062 0 1 -2081
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X7
timestamp 0
transform 1 0 6431 0 1 -2134
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X8
timestamp 0
transform 1 0 4586 0 1 -1869
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X9
timestamp 0
transform 1 0 4955 0 1 -1922
box -211 -420 211 420
use sky130_fd_pr__pfet_01v8_6FCS7L  X10
timestamp 0
transform 1 0 1634 0 1 -1436
box -211 -429 211 429
use sky130_fd_pr__pfet_01v8_ETRZ5W  X11
timestamp 0
transform 1 0 2003 0 1 -1489
box -211 -429 211 429
use sky130_fd_pr__pfet_01v8_6FCS7L  X12
timestamp 0
transform 1 0 158 0 1 -1224
box -211 -429 211 429
use sky130_fd_pr__pfet_01v8_ETRZ5W  X13
timestamp 0
transform 1 0 527 0 1 -1277
box -211 -429 211 429
use sky130_fd_pr__nfet_01v8_UJAU4L  X14
timestamp 0
transform 1 0 3848 0 1 -1763
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X15
timestamp 0
transform 1 0 4217 0 1 -1816
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_UJAU4L  X16
timestamp 0
transform 1 0 3110 0 1 -1657
box -211 -420 211 420
use sky130_fd_pr__nfet_01v8_44W2XU  X17
timestamp 0
transform 1 0 3479 0 1 -1710
box -211 -420 211 420
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 INN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 INP
port 4 nsew
<< end >>
